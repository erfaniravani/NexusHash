`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/19/2021 05:35:28 AM
// Design Name: 
// Module Name: test_bench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test_bench();

    reg clk;
    //reg [7:0] d;
    reg [1087:0] key;
    reg [1023:0] message;
    //reg [191:0] tweak;
    //reg [21503:0] subkey;
    wire [1023:0] oup;
    wire [63:0] mozp;
    wire [63:0] nonce;
    wire correct;
    //wire [1023:0] done;
    //wire [1087:0] key;
    connector CNCTR(clk,key,message,oup,mozp,nonce,correct);
    
    initial begin
        clk = 0;
        message = 1024'h0b87c738f85418020aeb2dc8f705eaf32f497e4eb506aacad70a51eb6b1db311da1c1342f2652ff2e29f01df55a6ddd340f30914dac10e3105476f7aa3989fc600000002010082667b04aa8a003dc787000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        //d = 8'd7;
        //#102
        //tweak = 192'h03000D02400008FF00000020870000FF000310A0000008;
        //subkey = 21504'd1900997572;
        key = 1088'h24b9d5b04edfc22ac530df071015100fbaa2d6bb0ca3b08207878b1fafa4cef774b7d109268e689380f5da9663621229967afe4d9a6387527d429271833937f0a39995d0acc6537ea3fc0a2e08a9aab2a0fd444162347c347a6494fa5c37c487b8b703a467f844161b0673fbea904d3cb68830dbc2a97498f1238495700021a22865eeb151832e72;
        //#4
        //subkey = 21504'd6854364338985098654;
        //key = 1088'h1B7A4E6E0DFDA99ACDE136B4D772C807690A1C1145FE576620BA18BF10E2584B89C2BDE3EC22AEC7FC44BA6825810316C823D73E9D71B706B12114950878B9B6CA7CE3B8ACA974A4502F5FD5522B7388DB8A6EF98F3D9DADD71E1132B95D485C2E248DC470E5E342365F98A64502119A89B5D42022CE0C702948DDB1FE45968BE8BB3254A7E2227A;
        //#4
        //subkey = 21504'd753087543136;
        //message = 1024'hBD1DD3D31E6BA2699655072155D642E0F17A80CEB86EB594FF5649866BFD457A64C940C6E197128C48971E4AAB73848BC19848A8326323E66E339FE3F81454B8B032AD1453302AEF8EC248370CE833B3E6C15AD2D93BA13758C25DB0F9AACFD9AEB301322D1E8A57046A8A28295AE7D18080FD19D3214BD21B926841B6E8B5FF;
        //#4
        //subkey = 21504'd1900997572;
        //message = 1024'hAB0CAEC403DA0B2E6DCE92682DE6770843A0F4803D406C35DD05BDD04553FFDBA51264C74D09926043BFAC6DA4A6CF6FDCE1AF1D7D0A2DEB5B2405D00F9449FA00000002019BFC7C7B03DE50003D9702000000000000031C00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        //#4
        //subkey = 21504'd6854364338985098654;
        //message = 1024'h40239A391A6507F87420CE999680C868BB2052B2E53194E167FD3DB5E9F4F55827D944C639253C84DA93129425AC3DFA3E08C20864EAA63670D12DD86264DCE400000002DB4B1BD67B0CF7DF003DA33F000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        //#4
        //subkey = 21504'd753087543136;
        //message = 1024'hBD1DD3D31E6BA2699655072155D642E0F17A80CEB86EB594FF5649866BFD457A64C940C6E197128C48971E4AAB73848BC19848A8326323E66E339FE3F81454B8B032AD1453302AEF8EC248370CE833B3E6C15AD2D93BA13758C25DB0F9AACFD9AEB301322D1E8A57046A8A28295AE7D18080FD19D3214BD21B926841B6E8B5FF;
        //#4
        //subkey = 21504'd1900997572;
        //message = 1024'b0;
        #2000 $stop;
    end
    
    always
    begin
        #2 clk = ~clk;
    end

endmodule
